module controller(
);

endmodule