module upcount2(
	input logic CLR, CLKb,
	output logic [1:0] CNT
);

endmodule