module ALU(
	input logic [9:0] OP,
	input logic [3:0] FN,
	input logic Ain, Gin, Gout, CLKb,
	output logic [9:0] Q
);

endmodule